///////////////////////////////////////////////////////////////////////////////////
///                                                                             /// 
///                      Events to APB Transaction Module                       ///
///                                                                             ///
///////////////////////////////////////////////////////////////////////////////////
///  This design detects a 3 bit overlapping serial palindrome sequence         ///
///                                                                             ///
///  Copyright 2025 Ujval Madhu, All rights reserved                            ///
///////////////////////////////////////////////////////////////////////////////////
//  CVS Log
//
//  Id: events_to_APB.v, v 1.0
//
//  $Date: 2024-02-05
//  $Revision: 1.0 $
//  $Author:  Ujval Madhu

module palindrome3b (
  input   logic        clk,
  input   logic        reset,

  input   logic        x_i,

  output  logic        palindrome_o
);


    
endmodule