///////////////////////////////////////////////////////////////////////////////////
///                                  ///
///                                                                             ///
///////////////////////////////////////////////////////////////////////////////////
///    Module:                                                               ///
///                                                                             ///
///   Copyright 2025 Ujval Madhu, All rights reserved                           ///
///////////////////////////////////////////////////////////////////////////////////
//  CVS Log
//
//  Id:  v 1.0
//
//  $Date: 2024-07-03
//  $Revision: 1.0 $
//  $Author:  Ujval Madhu

