///////////////////////////////////////////////////////////////////////////////////
///                                                                             ///
///              Testbench for 36-Bit Braun Multiplier                        ///
///                                                                             ///
///////////////////////////////////////////////////////////////////////////////////
///   Testbench Module: Verification using Randomized Stimulus,                 ///
///                     Functional Equivalence and Immediate Assertion          ///
///            This code is Generated by a Perl Script.                         ///
///                                                                             ///
///   Copyright (C) 2025 Ujval Madhu,                                           ///
///   This program is free software: you can redistribute it and/or modify      ///
///   it under the terms of the GNU General Public License as published by      ///
///   the Free Software Foundation, either version 3 of the License, or         ///
///   (at your option) any later version.                                       ///
///                                                                             ///
///   This program is distributed in the hope that it will be useful,           ///
///   but WITHOUT ANY WARRANTY; without even the implied warranty of            ///
///   MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the             ///
///   GNU General Public License for more details.                              ///
///                                                                             ///
///   You should have received a copy of the GNU General Public License         ///
///   along with this program.  If not, see <https://www.gnu.org/licenses/>.    ///
///                                                                             ///
///////////////////////////////////////////////////////////////////////////////////
//  CVS Log
//
//  Id: testbench.sv, v 1.0
//
//  $Date: 2025-4-7
//  $Revision: 1.0 
//  $Author:  Ujval Madhu


module testbench;

    parameter num_bits = 18;
    parameter num_tests = 100;

    reg [num_bits -1:0] in_a;
    reg [num_bits -1:0] in_b;
    
    reg [(2*num_bits) -1:0] prod;
    reg [(2*num_bits) -1:0] expected_prod;

    integer seed;

    // Instantiating the Braun Multiplier
    braun_mult bmx(.a(in_a), .b(in_b), .prod(prod));
    
    ////////////////////////////////
    //    Random Stimulus Test    //
    ////////////////////////////////

    initial begin
        seed = $urandom;
        $urandom(seed);              // Icarus doesn't support $srandom yet

        in_b = 18'b0;
        in_a = 18'b0;
        #10;
        
        for(int i = 1; i <= num_tests; i++) begin
            in_a = $urandom % (2**18 - 1);
            in_b = $urandom % (2**18 - 1);

            #10;

            $display("\n Random Test %0d", i);
            $display("Braun Multiplier Result: Input A: %d, Input B: %d, Product: %d", in_a, in_b, prod);

           //////////////////////// 
           // Functional Testing //
           ////////////////////////

            expected_prod =  in_a * in_b;

            assert(expected_prod == prod)
            else begin
                $error("Product Check Assertion error: Expected Product = %0d, but Obtained Product = %0d at %0t", expected_prod, prod, $time);
                $fatal;
            end
            
            #10;

        end

        $display("\nAll %0d Test cases Passed !!\n", num_tests);

    end

    // Generating Waveform Files
    initial begin
        $dumpfile("testbench.vcd");
        $dumpvars(0, testbench);
    end

endmodule
